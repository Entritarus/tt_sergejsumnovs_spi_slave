library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package data_types is
  alias sl is std_logic;
  alias slv is std_logic_vector;
  type aslv is array(integer range <>) of std_logic_vector;
end package data_types;

package body data_types is
end package body;
