/*
 * Copyright (c) 2025 Sergejs Umnovs
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_sergejsumnovs_spi_slave (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  test_component(clk, rst_n, uo_out);
  // All output pins must be assigned. If not used, assign to 0.
  assign uio_out = 0;
  assign uio_oe  = 0;

  //assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, ui_in, uio_in, uio_out, uio_oe, 1'b0};

  

endmodule
